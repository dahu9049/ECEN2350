module hexEncode(input [3:0] bin, output reg [7:0] hex);
    always @(bin) begin
        case(bin)
            4'b0000 : hex = 8'b11000000; // 0
            4'b0001 : hex = 8'b11111001; // 1
            4'b0010 : hex = 8'b10100100; // 2
            4'b0011 : hex = 8'b10110000; // 3
            4'b0100 : hex = 8'b10011001; // 4
            4'b0101 : hex = 8'b10010010; // 5
            4'b0110 : hex = 8'b10000010; // 6 
            4'b0111 : hex = 8'b11111000; // 7
            4'b1000 : hex = 8'b10000000; // 8
            4'b1001 : hex = 8'b10010000; // 9
            4'b1010 : hex = 8'b10001000; // 10
            4'b1011 : hex = 8'b10000011; // 11
            4'b1100 : hex = 8'b11000110; // 12
            4'b1101 : hex = 8'b10100001; // 13
            4'b1110 : hex = 8'b10000110; // 14
            4'b1111 : hex = 8'b10001110; // 15
        endcase
    end
endmodule